**.subckt tb_inverter vin vout
*.opin vin
*.opin vout
x1 net1 vin vout GND inverter
V1 net1 GND 1.8
V2 vin GND PWL(0 0 20n 0 900n 1.8)
**** begin user architecture code

.lib /usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 1n 1u
plot V(vout) V(vin)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
* sym_path: /home/shabbarvejlani/workshop/inverter/xschem/inverter.sym
* sch_path: /home/shabbarvejlani/workshop/inverter/xschem/inverter.sch
.subckt inverter  vdd vin vout vss
*.ipin vin
*.iopin vdd
*.iopin vss
*.opin vout
XM3 vout vin vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=4.5 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

.GLOBAL GND
** flattened .save nodes
.end
